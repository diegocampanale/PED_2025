module distributore();

endmodule